** test circuit for selector
.include General model.cir
* Use this for repeating pulses


.param vread = 0.08
.param vset = 1
.param tdelay = 1ms
.param tedge = 1us
.param ton = 1ms
.param ttotal = 10ms
.param cycles = 1
* selector
*Syntax: Vxxx n+ n- PULSE(V1 V2 Tdelay Trise Tfall Ton Tperiod Ncycles)
V1 p 0 pulse({vread} {vset} 1ms {tedge} {tedge} {ton} {ttotal} {cycles})
XSelector p 0 memristor n = 2, m=2, h1= 10e-9, h2 =5e-9, alpha=3.589e-12, beta=2.659e-12, sigma=1.061e-8, eta = 1.25e-16, theta = 0.32, Ron = 8.6e3, Roff = 1e9, cc = 100e-6

* Transient simulation
* Transient simulation
.TRAN 1us {ttotal*cycles} 0 .0001ms
.PROBE
.END





