* Diffusive memristor test: multiple voltage pulses input

* Model parameters
.param alpha=0.1
.param lamda=0.1
.param Ron=1.7e4
.param Roff=1e10
.param mu=16
.param beta=0.2
.param gamma1=50
.param gamma2=0.42
.param eta=0.01

* Optional noise controls
.param dt=1e-3
.param kappa=200
.param m=2
.param eps=1e-12

* Multi-pulse voltage stimulus
.param Vamp=0.8
.param tdelay=1ms
.param trise=10us
.param tfall=10us
.param ton=0.8s
.param tperiod=1.1s
.param cycles=30
.param tstop={tdelay + cycles*tperiod + 10ms}

.include "Diffusive_model_core.cir"

Vin in 0 PULSE(0 {Vamp} {tdelay} {trise} {tfall} {ton} {tperiod} {cycles})
Rs in p 50
Rp p n 1e7
Cp2 p n 1e-6
Vgnd n 0 0

.tran 0 {tstop} 0 0.1ms

* Save both input pulse and device response
.save V(in) I(Vin) V(p) V(n) V(f) V(r) I(BIMx)
.plot tran V(in) I(Vin) V(p) V(f) V(r) I(BIMx)
.probe
.end
