** Selector model
.subckt memristor p minus
* Selector model UMass Threshold Switching Device
* Ye, IEDM Lab/Yang group, UMass Amherst, 2019
* p & n are the terminals, Selector is the device name


*** If you want a faster/low threshold voltage, you can increase down alpha and eta, or decrease beta and theta.  Also h1, h2 will afftect the turn-on and turn-off voltage.

*** if you need to change to non-linearity of conductance, you can change the h_lambda.


**  h0 is the initial length, hmax is the max length
**  h1 is the turn on length, h2 is the turn off length
**  n, h_lambda are the exponetial parameters
**  alpha, beta are the pre-exponetial parameters
.param n = {n}
.param h0 = 0
.param hmax = 15e-9
.param h1 = {h1}
.param h2 = {h2}
.param h_lambda = 1e-8
.param alpha = {alpha}
.param beta = {beta}

**  s0 is the initial length,
**  h1 is the turn on length,
**  m is the exponetial parameters
**  eta, theta are the pre-exponetial parameters
.param m = {m}
.param s0 = 1e-16
.param smin = 0.9999*s0
.param smax = 1.001*s0
.param sigma = {sigma}
.param eta = {eta}
.param theta = {theta}

** Ron, Roff are the on/off resistance
.param Ron = 8.6e3
.param Roff = 1e9
* current compliance
.param cc = 100e-6

*** Dynamic equation. How the state variable h/s will change given external stimulus.
Gh 0 h_ value= {dhdt(V(p), V(h), V(s_))}
Ch h_ 0 1 IC={0}
Rh h h_ 0.000000000001
Eh h 0 value = {limit(V(h_), -1e-11, 1.0001*hmax)}

Gs 0 s_ value= {dsdt(V(p), V(h), V(s))}
Cs s_ 0 1 IC={s0}
Rs s s_ 0.000000000001
Es s 0 value = {limit(V(s_), smin, smax)}


** dhdt_, dsdt_, the switching conditions
.func dhdt(v, h, s) {if(iout(v, h, s)< cc, dhdt_(v, h, s), 0)}
.func dsdt(v, h, s) {dsdt_(v, h, s)}

.func dhdt_(v, h, s) {if(h<hmax | (h>=hmax & dsdt__(v, h, s)<0 & s <= s0) , dhdt__(v, h, s), 0)}
.func dsdt_(v, h, s) {if(h<hmax | (h>=hmax & dsdt__(v, h, s)<0 & s <= s0) , 0, dsdt__(v, h, s))}


** dhdt, dsdt. the swtiching rate of h, s
.func dhdt__(v, h, s) {alpha*pow(v, n)*1/(sqrt(2*Pi)*sigma)*exp(-1/2*pow((h-h1)/sigma, 2))-beta*h/hmax*1/(sqrt(2*Pi)*sigma)*exp(-1/2*pow((h-h2)/sigma, 2))}
.func dsdt__(v, h, s) {eta*pow(v, m)*exp(-s)-theta*s}

** memristance. the definition of the memristance
.func memristance(h, s) {Ron*h/hmax * sqrt(s0/s) + Roff*(exp(hmax/h_lambda-h/h_lambda)-1)/(exp(hmax/h_lambda)-1)}

.func iout(v, h, s) = min(v/memristance(limit(h,0, hmax), limit(s, smin, smax)), cc)
***  the output current between p, 0.
*BIMx plus minus I = dhdt_(V(p, n), V(h), V(s))
BIx p minus I = iout(V(p)-V(minus), v(h), v(s))
.ends




