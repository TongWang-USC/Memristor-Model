** test circuit for selector
.include General model.cir
* Use this for repeating pulses


.param vread = 0.1
.param vset = 2
.param vreset = -2
.param tdelay = 100us
.param tedge = 1us
.param ton = 50us
.param ttotal = 0.5ms
.param cycles = 2
* memristor
*Syntax: Vxxx n+ n- PULSE(V1 V2 Tdelay Trise Tfall Ton Tperiod Ncycles)
V1 p p1 pulse(0 {vset-vread} {tdelay} {tedge} {tedge} {ton} {ttotal} {cycles})
V2 p1 p2 pulse(0 {vreset-vread} {2*tdelay+2*tedge+ton} {tedge} {tedge} {ton} {ttotal} {cycles})
V3 p2 0 pulse(0 {vread} 0us {tedge} {tedge} 15ms {ttotal} {cycles})


XBipolar p 0 memristor n = 3, m = 5, h1 = 1e-9, h2=5e-9, alpha=1.329e-11, beta=2.659e-13, sigma=1.061e-08, eta = 1.25e-16, theta = 0.32, Ron = 0.47e3, Roff = 1.7e3, cc = 1e-2

* Transient simulation
* Transient simulation
.TRAN 1us {ttotal*cycles} 0 .0001ms
.PROBE
.END





